

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

-- Sine lookup table. Input is 0 to 2^24-1 => 0 to 2pi
-- Output is -2^23 to 2^23-1 => -1 to ~1
entity sine_lookup is
  port (
    counter_i : in unsigned(7 downto 0);
    freq_o : out std_logic_vector(23 downto 0)
    );
end entity;

architecture rtl of sine_lookup is

  type LUT_t is array (256 downto 0) of signed(23 downto 0);

  signal LUT : LUT_t;

begin

    freq_o <= std_logic_vector(LUT(to_integer(unsigned(counter_i))));

    LUT(0) <= to_signed(0, 24);
    LUT(1) <= to_signed(205866, 24);
    LUT(2) <= to_signed(411609, 24);
    LUT(3) <= to_signed(617104, 24);
    LUT(4) <= to_signed(822227, 24);
    LUT(5) <= to_signed(1026855, 24);
    LUT(6) <= to_signed(1230864, 24);
    LUT(7) <= to_signed(1434132, 24);
    LUT(8) <= to_signed(1636536, 24);
    LUT(9) <= to_signed(1837954, 24);
    LUT(10) <= to_signed(2038265, 24);
    LUT(11) <= to_signed(2237348, 24);
    LUT(12) <= to_signed(2435084, 24);
    LUT(13) <= to_signed(2631353, 24);
    LUT(14) <= to_signed(2826036, 24);
    LUT(15) <= to_signed(3019018, 24);
    LUT(16) <= to_signed(3210181, 24);
    LUT(17) <= to_signed(3399410, 24);
    LUT(18) <= to_signed(3586592, 24);
    LUT(19) <= to_signed(3771613, 24);
    LUT(20) <= to_signed(3954362, 24);
    LUT(21) <= to_signed(4134729, 24);
    LUT(22) <= to_signed(4312606, 24);
    LUT(23) <= to_signed(4487885, 24);
    LUT(24) <= to_signed(4660460, 24);
    LUT(25) <= to_signed(4830229, 24);
    LUT(26) <= to_signed(4997087, 24);
    LUT(27) <= to_signed(5160936, 24);
    LUT(28) <= to_signed(5321676, 24);
    LUT(29) <= to_signed(5479210, 24);
    LUT(30) <= to_signed(5633444, 24);
    LUT(31) <= to_signed(5784285, 24);
    LUT(32) <= to_signed(5931641, 24);
    LUT(33) <= to_signed(6075424, 24);
    LUT(34) <= to_signed(6215548, 24);
    LUT(35) <= to_signed(6351928, 24);
    LUT(36) <= to_signed(6484481, 24);
    LUT(37) <= to_signed(6613129, 24);
    LUT(38) <= to_signed(6737793, 24);
    LUT(39) <= to_signed(6858398, 24);
    LUT(40) <= to_signed(6974872, 24);
    LUT(41) <= to_signed(7087145, 24);
    LUT(42) <= to_signed(7195149, 24);
    LUT(43) <= to_signed(7298818, 24);
    LUT(44) <= to_signed(7398091, 24);
    LUT(45) <= to_signed(7492908, 24);
    LUT(46) <= to_signed(7583211, 24);
    LUT(47) <= to_signed(7668947, 24);
    LUT(48) <= to_signed(7750063, 24);
    LUT(49) <= to_signed(7826510, 24);
    LUT(50) <= to_signed(7898244, 24);
    LUT(51) <= to_signed(7965219, 24);
    LUT(52) <= to_signed(8027397, 24);
    LUT(53) <= to_signed(8084739, 24);
    LUT(54) <= to_signed(8137211, 24);
    LUT(55) <= to_signed(8184782, 24);
    LUT(56) <= to_signed(8227423, 24);
    LUT(57) <= to_signed(8265107, 24);
    LUT(58) <= to_signed(8297813, 24);
    LUT(59) <= to_signed(8325521, 24);
    LUT(60) <= to_signed(8348214, 24);
    LUT(61) <= to_signed(8365878, 24);
    LUT(62) <= to_signed(8378503, 24);
    LUT(63) <= to_signed(8386081, 24);
    LUT(64) <= to_signed(8388608, 24);
    LUT(65) <= to_signed(8386081, 24);
    LUT(66) <= to_signed(8378503, 24);
    LUT(67) <= to_signed(8365878, 24);
    LUT(68) <= to_signed(8348214, 24);
    LUT(69) <= to_signed(8325521, 24);
    LUT(70) <= to_signed(8297813, 24);
    LUT(71) <= to_signed(8265107, 24);
    LUT(72) <= to_signed(8227423, 24);
    LUT(73) <= to_signed(8184782, 24);
    LUT(74) <= to_signed(8137211, 24);
    LUT(75) <= to_signed(8084739, 24);
    LUT(76) <= to_signed(8027397, 24);
    LUT(77) <= to_signed(7965219, 24);
    LUT(78) <= to_signed(7898244, 24);
    LUT(79) <= to_signed(7826510, 24);
    LUT(80) <= to_signed(7750063, 24);
    LUT(81) <= to_signed(7668947, 24);
    LUT(82) <= to_signed(7583211, 24);
    LUT(83) <= to_signed(7492908, 24);
    LUT(84) <= to_signed(7398091, 24);
    LUT(85) <= to_signed(7298818, 24);
    LUT(86) <= to_signed(7195149, 24);
    LUT(87) <= to_signed(7087145, 24);
    LUT(88) <= to_signed(6974872, 24);
    LUT(89) <= to_signed(6858398, 24);
    LUT(90) <= to_signed(6737793, 24);
    LUT(91) <= to_signed(6613129, 24);
    LUT(92) <= to_signed(6484481, 24);
    LUT(93) <= to_signed(6351928, 24);
    LUT(94) <= to_signed(6215548, 24);
    LUT(95) <= to_signed(6075424, 24);
    LUT(96) <= to_signed(5931641, 24);
    LUT(97) <= to_signed(5784285, 24);
    LUT(98) <= to_signed(5633444, 24);
    LUT(99) <= to_signed(5479210, 24);
    LUT(100) <= to_signed(5321676, 24);
    LUT(101) <= to_signed(5160936, 24);
    LUT(102) <= to_signed(4997087, 24);
    LUT(103) <= to_signed(4830229, 24);
    LUT(104) <= to_signed(4660460, 24);
    LUT(105) <= to_signed(4487885, 24);
    LUT(106) <= to_signed(4312606, 24);
    LUT(107) <= to_signed(4134729, 24);
    LUT(108) <= to_signed(3954362, 24);
    LUT(109) <= to_signed(3771613, 24);
    LUT(110) <= to_signed(3586592, 24);
    LUT(111) <= to_signed(3399410, 24);
    LUT(112) <= to_signed(3210181, 24);
    LUT(113) <= to_signed(3019018, 24);
    LUT(114) <= to_signed(2826036, 24);
    LUT(115) <= to_signed(2631353, 24);
    LUT(116) <= to_signed(2435084, 24);
    LUT(117) <= to_signed(2237348, 24);
    LUT(118) <= to_signed(2038265, 24);
    LUT(119) <= to_signed(1837954, 24);
    LUT(120) <= to_signed(1636536, 24);
    LUT(121) <= to_signed(1434132, 24);
    LUT(122) <= to_signed(1230864, 24);
    LUT(123) <= to_signed(1026855, 24);
    LUT(124) <= to_signed(822227, 24);
    LUT(125) <= to_signed(617104, 24);
    LUT(126) <= to_signed(411609, 24);
    LUT(127) <= to_signed(205866, 24);
    LUT(128) <= to_signed(0, 24);
    LUT(129) <= to_signed(-205866, 24);
    LUT(130) <= to_signed(-411609, 24);
    LUT(131) <= to_signed(-617104, 24);
    LUT(132) <= to_signed(-822227, 24);
    LUT(133) <= to_signed(-1026855, 24);
    LUT(134) <= to_signed(-1230864, 24);
    LUT(135) <= to_signed(-1434132, 24);
    LUT(136) <= to_signed(-1636536, 24);
    LUT(137) <= to_signed(-1837954, 24);
    LUT(138) <= to_signed(-2038265, 24);
    LUT(139) <= to_signed(-2237348, 24);
    LUT(140) <= to_signed(-2435084, 24);
    LUT(141) <= to_signed(-2631353, 24);
    LUT(142) <= to_signed(-2826036, 24);
    LUT(143) <= to_signed(-3019018, 24);
    LUT(144) <= to_signed(-3210181, 24);
    LUT(145) <= to_signed(-3399410, 24);
    LUT(146) <= to_signed(-3586592, 24);
    LUT(147) <= to_signed(-3771613, 24);
    LUT(148) <= to_signed(-3954362, 24);
    LUT(149) <= to_signed(-4134729, 24);
    LUT(150) <= to_signed(-4312606, 24);
    LUT(151) <= to_signed(-4487885, 24);
    LUT(152) <= to_signed(-4660460, 24);
    LUT(153) <= to_signed(-4830229, 24);
    LUT(154) <= to_signed(-4997087, 24);
    LUT(155) <= to_signed(-5160936, 24);
    LUT(156) <= to_signed(-5321676, 24);
    LUT(157) <= to_signed(-5479210, 24);
    LUT(158) <= to_signed(-5633444, 24);
    LUT(159) <= to_signed(-5784285, 24);
    LUT(160) <= to_signed(-5931641, 24);
    LUT(161) <= to_signed(-6075424, 24);
    LUT(162) <= to_signed(-6215548, 24);
    LUT(163) <= to_signed(-6351928, 24);
    LUT(164) <= to_signed(-6484481, 24);
    LUT(165) <= to_signed(-6613129, 24);
    LUT(166) <= to_signed(-6737793, 24);
    LUT(167) <= to_signed(-6858398, 24);
    LUT(168) <= to_signed(-6974872, 24);
    LUT(169) <= to_signed(-7087145, 24);
    LUT(170) <= to_signed(-7195149, 24);
    LUT(171) <= to_signed(-7298818, 24);
    LUT(172) <= to_signed(-7398091, 24);
    LUT(173) <= to_signed(-7492908, 24);
    LUT(174) <= to_signed(-7583211, 24);
    LUT(175) <= to_signed(-7668947, 24);
    LUT(176) <= to_signed(-7750063, 24);
    LUT(177) <= to_signed(-7826510, 24);
    LUT(178) <= to_signed(-7898244, 24);
    LUT(179) <= to_signed(-7965219, 24);
    LUT(180) <= to_signed(-8027397, 24);
    LUT(181) <= to_signed(-8084739, 24);
    LUT(182) <= to_signed(-8137211, 24);
    LUT(183) <= to_signed(-8184782, 24);
    LUT(184) <= to_signed(-8227423, 24);
    LUT(185) <= to_signed(-8265107, 24);
    LUT(186) <= to_signed(-8297813, 24);
    LUT(187) <= to_signed(-8325521, 24);
    LUT(188) <= to_signed(-8348214, 24);
    LUT(189) <= to_signed(-8365878, 24);
    LUT(190) <= to_signed(-8378503, 24);
    LUT(191) <= to_signed(-8386081, 24);
    LUT(192) <= to_signed(-8388608, 24);
    LUT(193) <= to_signed(-8386081, 24);
    LUT(194) <= to_signed(-8378503, 24);
    LUT(195) <= to_signed(-8365878, 24);
    LUT(196) <= to_signed(-8348214, 24);
    LUT(197) <= to_signed(-8325521, 24);
    LUT(198) <= to_signed(-8297813, 24);
    LUT(199) <= to_signed(-8265107, 24);
    LUT(200) <= to_signed(-8227423, 24);
    LUT(201) <= to_signed(-8184782, 24);
    LUT(202) <= to_signed(-8137211, 24);
    LUT(203) <= to_signed(-8084739, 24);
    LUT(204) <= to_signed(-8027397, 24);
    LUT(205) <= to_signed(-7965219, 24);
    LUT(206) <= to_signed(-7898244, 24);
    LUT(207) <= to_signed(-7826510, 24);
    LUT(208) <= to_signed(-7750063, 24);
    LUT(209) <= to_signed(-7668947, 24);
    LUT(210) <= to_signed(-7583211, 24);
    LUT(211) <= to_signed(-7492908, 24);
    LUT(212) <= to_signed(-7398091, 24);
    LUT(213) <= to_signed(-7298818, 24);
    LUT(214) <= to_signed(-7195149, 24);
    LUT(215) <= to_signed(-7087145, 24);
    LUT(216) <= to_signed(-6974872, 24);
    LUT(217) <= to_signed(-6858398, 24);
    LUT(218) <= to_signed(-6737793, 24);
    LUT(219) <= to_signed(-6613129, 24);
    LUT(220) <= to_signed(-6484481, 24);
    LUT(221) <= to_signed(-6351928, 24);
    LUT(222) <= to_signed(-6215548, 24);
    LUT(223) <= to_signed(-6075424, 24);
    LUT(224) <= to_signed(-5931641, 24);
    LUT(225) <= to_signed(-5784285, 24);
    LUT(226) <= to_signed(-5633444, 24);
    LUT(227) <= to_signed(-5479210, 24);
    LUT(228) <= to_signed(-5321676, 24);
    LUT(229) <= to_signed(-5160936, 24);
    LUT(230) <= to_signed(-4997087, 24);
    LUT(231) <= to_signed(-4830229, 24);
    LUT(232) <= to_signed(-4660460, 24);
    LUT(233) <= to_signed(-4487885, 24);
    LUT(234) <= to_signed(-4312606, 24);
    LUT(235) <= to_signed(-4134729, 24);
    LUT(236) <= to_signed(-3954362, 24);
    LUT(237) <= to_signed(-3771613, 24);
    LUT(238) <= to_signed(-3586592, 24);
    LUT(239) <= to_signed(-3399410, 24);
    LUT(240) <= to_signed(-3210181, 24);
    LUT(241) <= to_signed(-3019018, 24);
    LUT(242) <= to_signed(-2826036, 24);
    LUT(243) <= to_signed(-2631353, 24);
    LUT(244) <= to_signed(-2435084, 24);
    LUT(245) <= to_signed(-2237348, 24);
    LUT(246) <= to_signed(-2038265, 24);
    LUT(247) <= to_signed(-1837954, 24);
    LUT(248) <= to_signed(-1636536, 24);
    LUT(249) <= to_signed(-1434132, 24);
    LUT(250) <= to_signed(-1230864, 24);
    LUT(251) <= to_signed(-1026855, 24);
    LUT(252) <= to_signed(-822227, 24);
    LUT(253) <= to_signed(-617104, 24);
    LUT(254) <= to_signed(-411609, 24);
    LUT(255) <= to_signed(-205866, 24);
end rtl;
